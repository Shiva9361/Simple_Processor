module set_less_then(input a,input b);
endmodule